*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TB_JNW_GR03_AMP_lpe.spi
#else
.include ../../../work/xsch/TB_JNW_GR03_AMP.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}
.param mc_mm_switch=0
.param mc_pr_switch=0

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
*.save all
.save v(out_amp)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0
op

ac dec 50 1 1e9

let vo_mag = db(v(out_amp))
write {cicname}.raw
quit
.endc
.end
