*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_GR03_lpe.spi
#else
.include ../../../work/xsch/JNW_GR03.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  VSS   dc 1.8
VRST RST  0     pulse(0 1.8 0 2n 2n 1u 10u 1) 
VCLK  CLK 0     pulse(0 1.8 5n 1n 1n 6n 20n)


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi
.include ../svinst.spi
*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

.save v(OUT)
.save v(RST_CAP)
.save v(COMP)


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0



set fend = .raw
* foreach vtemp -25 0 25 50 75 100 120
foreach vtemp -25 50 120
    option temp=$vtemp
    tran 1n 10u 1n
    write {cicname}_$vtemp$fend
end

quit
.endc
.end
