magic
tech sky130A
magscale 1 2
timestamp 1744301330
<< error_p >>
rect 12177 13192 12930 13250
<< error_s >>
rect 8484 19560 8536 20616
rect 10749 20214 10755 20220
rect 10743 20208 10749 20214
rect 10743 20150 10749 20156
rect 10749 20144 10755 20150
rect 11929 20124 12179 20932
rect 12273 20214 12279 20220
rect 12267 20208 12273 20214
rect 12267 20150 12273 20156
rect 12273 20144 12279 20150
rect 13455 20124 13703 20932
rect 13799 20214 13805 20220
rect 13793 20208 13799 20214
rect 13793 20150 13799 20156
rect 13799 20144 13805 20150
rect 14980 20128 15229 20936
rect 19131 20884 19264 20890
rect 19170 20830 19210 20836
rect 19170 20796 19176 20802
rect 15324 20218 15330 20224
rect 15318 20212 15324 20218
rect 18088 20172 18094 20178
rect 18082 20166 18088 20172
rect 15318 20154 15324 20160
rect 15324 20148 15330 20154
rect 14726 20124 14975 20128
rect 10405 19876 11925 20124
rect 11929 19876 13449 20124
rect 13455 19876 14975 20124
rect 14980 19880 16500 20128
rect 18082 20108 18088 20114
rect 18088 20102 18094 20108
rect 11929 18814 12179 19870
rect 12273 18924 12279 18930
rect 12267 18918 12273 18924
rect 12267 18860 12273 18866
rect 12273 18854 12279 18860
rect 13455 18814 13703 19870
rect 14862 18916 14868 18922
rect 14856 18910 14862 18916
rect 14980 18818 15229 19874
rect 17744 19834 19264 20082
rect 19385 20076 19518 20884
rect 19729 20166 19735 20172
rect 19723 20160 19729 20166
rect 19723 20102 19729 20108
rect 19729 20096 19735 20102
rect 20909 20076 21159 20884
rect 21253 20166 21259 20172
rect 21247 20160 21253 20166
rect 21247 20102 21253 20108
rect 21253 20096 21259 20102
rect 22435 20076 22683 20884
rect 22779 20166 22785 20172
rect 22773 20160 22779 20166
rect 22773 20102 22779 20108
rect 22779 20096 22785 20102
rect 19385 19828 20905 20076
rect 20909 19828 22429 20076
rect 22435 19828 23955 20076
rect 19131 19822 19264 19828
rect 19385 18772 19518 19822
rect 20909 19484 21159 19822
rect 20909 18766 21056 19484
rect 22435 18766 22683 19822
rect 12019 16772 12021 16776
rect 13545 16772 13547 16776
rect 11985 16738 12021 16742
rect 13511 16738 13547 16742
rect 10885 16570 11065 16736
rect 12409 16570 12589 16736
rect 13935 16570 14115 16736
rect 10883 16556 11065 16570
rect 12407 16556 12589 16570
rect 13933 16556 14115 16570
rect 15460 16564 15640 16740
rect 20999 16724 21001 16728
rect 22525 16724 22527 16728
rect 20965 16690 21001 16694
rect 22491 16690 22527 16694
rect 15460 16560 15663 16564
rect 10883 16390 11063 16556
rect 12407 16390 12587 16556
rect 13933 16390 14113 16556
rect 11983 16384 12019 16388
rect 13509 16384 13545 16388
rect 15483 16384 15663 16560
rect 16583 16378 16619 16382
rect 18109 16378 18145 16382
rect 12017 16350 12019 16354
rect 13543 16350 13545 16354
rect 16617 16344 16619 16348
rect 18143 16344 18145 16348
rect 10403 13256 11923 13504
rect 11927 13256 12066 14312
rect 13453 13504 13701 14312
rect 14749 14306 14973 14312
rect 12177 13256 13447 13504
rect 13453 13256 14973 13504
rect 15003 13498 15227 14306
rect 16527 13498 16777 14306
rect 16871 14260 16877 14266
rect 16865 14254 16871 14260
rect 16865 14196 16871 14202
rect 16871 14190 16877 14196
rect 18053 13498 18301 14306
rect 15003 13250 16523 13498
rect 16527 13250 18047 13498
rect 18053 13250 19573 13498
rect 11927 13192 12066 13250
rect 10747 12976 10753 12982
rect 10741 12970 10747 12976
rect 10741 12912 10747 12918
rect 10747 12906 10753 12912
rect 11927 12194 12177 13192
rect 12271 12976 12277 12982
rect 12265 12970 12271 12976
rect 12265 12912 12271 12918
rect 12271 12906 12277 12912
rect 13453 12194 13701 13250
rect 14749 13244 14973 13250
rect 13797 12976 13803 12982
rect 13791 12970 13797 12976
rect 13791 12912 13797 12918
rect 13797 12906 13803 12912
rect 15003 12194 15227 13244
rect 15347 12970 15353 12976
rect 15341 12964 15347 12970
rect 15341 12906 15347 12912
rect 15347 12900 15353 12906
rect 15347 12356 15368 12364
rect 15319 12328 15340 12336
rect 16527 12188 16777 13244
rect 16871 12970 16877 12976
rect 16865 12964 16871 12970
rect 16865 12906 16871 12912
rect 16871 12900 16877 12906
rect 18053 12188 18301 13244
rect 18397 12970 18403 12976
rect 18391 12964 18397 12970
rect 18391 12906 18397 12912
rect 18397 12900 18403 12906
<< error_ps >>
rect 21056 18766 21159 19484
rect 21253 18876 21259 18882
rect 21247 18870 21253 18876
rect 21247 18812 21253 18818
rect 21253 18806 21259 18812
rect 12066 13256 12177 14312
rect 12271 14266 12277 14272
rect 12265 14260 12271 14266
rect 12265 14202 12271 14208
rect 12271 14196 12277 14202
rect 12066 13192 12177 13250
<< locali >>
rect 6850 20524 10638 21062
rect 14232 21022 16624 21070
rect 14232 20878 24470 21022
rect 16228 20830 24470 20878
rect 7822 18474 9894 18530
rect 7822 18338 10594 18474
rect 9686 17590 10594 18338
rect 10514 16424 16388 16698
rect 19416 15800 23844 16544
rect 24278 12288 24470 20830
rect 14480 12056 15814 12248
rect 19146 12096 24470 12288
<< metal1 >>
rect 10158 21158 16028 21350
rect 10158 19726 10350 21158
rect 15836 20528 16028 21158
rect 18600 20432 18792 21294
rect 23320 20520 23406 20584
rect 23470 20520 23476 20584
rect 8382 19524 8892 19588
rect 9342 19584 9406 19590
rect 7630 19248 7694 19254
rect 7630 19178 7694 19184
rect 8382 18194 8446 19524
rect 10158 19534 10822 19726
rect 9342 19514 9406 19520
rect 9406 11932 9470 18882
rect 14311 18724 14862 18916
rect 15054 18724 15386 18916
rect 15836 18696 18152 18888
rect 18600 18626 19796 18818
rect 23291 18644 23950 18836
rect 11514 17376 11520 17440
rect 11584 17376 11590 17440
rect 10170 16594 10362 16600
rect 10170 14442 10362 16402
rect 11520 16282 11584 17376
rect 11520 16212 11584 16218
rect 16490 16794 16554 16800
rect 16490 15920 16554 16730
rect 16490 15850 16554 15856
rect 18930 15078 18994 15084
rect 18930 14934 18994 15014
rect 10170 14250 10806 14442
rect 14309 14348 15406 14398
rect 14309 14284 14762 14348
rect 14826 14284 15406 14348
rect 14309 14206 15406 14284
rect 18934 12458 19042 12522
rect 19106 12458 19112 12522
rect 14744 12336 14808 12342
rect 14808 12272 15270 12336
rect 15334 12272 15340 12336
rect 14744 12266 14808 12272
rect 15272 11932 15336 11938
rect 9406 11868 15272 11932
rect 15272 11862 15336 11868
<< via1 >>
rect 23406 20520 23470 20584
rect 7630 19184 7694 19248
rect 9342 19520 9406 19584
rect 14862 18724 15054 18916
rect 11520 17376 11584 17440
rect 10170 16402 10362 16594
rect 11520 16218 11584 16282
rect 16490 16730 16554 16794
rect 16490 15856 16554 15920
rect 18930 15014 18994 15078
rect 14762 14284 14826 14348
rect 19042 12458 19106 12522
rect 14744 12272 14808 12336
rect 15270 12272 15334 12336
rect 15272 11868 15336 11932
<< metal2 >>
rect 18470 20744 23470 20808
rect 18470 20108 18534 20744
rect 23406 20584 23470 20744
rect 23406 20514 23470 20520
rect 9336 19520 9342 19584
rect 9406 19520 10276 19584
rect 7624 19184 7630 19248
rect 7694 19184 10058 19248
rect 9994 17112 10058 19184
rect 10212 17450 10276 19520
rect 10212 17386 10479 17450
rect 11520 17440 11584 17446
rect 11108 17376 11520 17440
rect 11520 17370 11584 17376
rect 9994 17048 10469 17112
rect 9994 15740 10058 17048
rect 14862 16594 15054 18724
rect 10164 16402 10170 16594
rect 10362 16402 15054 16594
rect 15710 16354 15774 17454
rect 18854 17338 19459 17402
rect 18854 16794 18918 17338
rect 16484 16730 16490 16794
rect 16554 16730 18918 16794
rect 15710 16290 19222 16354
rect 11514 16218 11520 16282
rect 11584 16218 15070 16282
rect 15006 16008 15070 16218
rect 14762 15856 16490 15920
rect 16554 15856 16560 15920
rect 9994 15676 10646 15740
rect 14762 14348 14826 15856
rect 14762 14278 14826 14284
rect 14190 12336 14254 12976
rect 14190 12272 14744 12336
rect 14808 12272 14814 12336
rect 15013 11796 15077 15734
rect 19158 15078 19222 16290
rect 18924 15014 18930 15078
rect 18994 15014 19222 15078
rect 19042 12522 19106 12528
rect 15270 12336 15334 12342
rect 19042 12336 19106 12458
rect 15334 12272 19106 12336
rect 15270 12266 15334 12272
rect 19385 11932 19449 17064
rect 15266 11868 15272 11932
rect 15336 11868 19449 11932
use JNW_GR03_NAND  x1 ../JNW_GR03_SKY130A
timestamp 1744282624
transform 1 0 14004 0 1 16836
box 976 -288 2500 4238
use JNW_GR03_NAND3  x2 ../JNW_GR03_SKY130A
timestamp 1744283476
transform 1 0 9269 0 1 16164
box 1107 374 5710 4910
use JNW_GR03_NAND3  x3
timestamp 1744283476
transform 1 0 9267 0 -1 16962
box 1107 374 5710 4910
use JNW_GR03_NAND3  x4
timestamp 1744283476
transform 1 0 13867 0 -1 16956
box 1107 374 5710 4910
use JNW_GR03_NAND3  x5
timestamp 1744283476
transform 1 0 18249 0 1 16116
box 1107 374 5710 4910
use JNW_GR03_NOT  x6 ../JNW_GR03_SKY130A
timestamp 1744281465
transform 0 -1 9876 1 0 18592
box -262 -128 2140 1392
use JNW_GR03_NOT  x7
timestamp 1744281465
transform 0 -1 8154 1 0 18592
box -262 -128 2140 1392
use JNW_GR03_NAND  x8
timestamp 1744282624
transform 1 0 16768 0 1 16790
box 976 -288 2500 4238
<< labels >>
flabel space 15012 11800 15062 12002 0 FreeSans 1600 0 0 0 D
port 0 nsew
flabel metal1 18600 21102 18792 21294 0 FreeSans 1600 0 0 0 Q
port 1 nsew
flabel metal1 23758 18644 23950 18836 0 FreeSans 1600 0 0 0 NOT_Q
port 2 nsew
flabel space 6844 20604 8346 21036 0 FreeSans 1600 0 0 0 VDD
port 3 nsew
flabel locali 9690 17698 9946 18446 0 FreeSans 1600 0 0 0 VSS
port 4 nsew
flabel space 7112 19374 7158 19790 0 FreeSans 1600 0 0 0 CLK
port 5 nsew
flabel metal1 8382 18194 8446 18258 0 FreeSans 1600 0 0 0 RST
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 69120 800
<< end >>
