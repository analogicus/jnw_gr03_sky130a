*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_GR03_AMP_lpe.spi
#else
.include ../../../work/xsch/JNW_GR03_AMP.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
* TNOM=27: Sets the nominal temperature to 27°C.
* GMIN=1e-15: Sets the minimum conductance to avoid floating nodes.
* reltol=1e-3: Sets the relative tolerance for iterative solutions.
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3


*-----------------------------------------------------------------
* PARAMETERS
* TRF = 10p: Defines a parameter for rise/fall time.
* AVDD: Defines a parameter for the supply voltage, which is set to {vdda}
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}   
* VDD_1V8 is the port name 
VIN  VIN  0     SIN(0 0.1 1k)  ; Input signal
VIP  VIP  0     dc 0 
*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save i(VDD) v(VIN) v(VIP) v(VO)


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 1n 10u
write
quit


.endc

.end
