magic
tech sky130A
magscale 1 2
timestamp 1744305162
<< metal1 >>
rect 9866 13834 9941 15787
rect 20298 13836 20365 15765
rect 30790 13862 30857 15845
rect 41310 13864 41377 15835
rect 8025 13767 9941 13834
rect 18476 13769 20365 13836
rect 29009 13795 30857 13862
rect 39466 13797 41377 13864
rect 51772 13862 51839 15835
rect 62260 13864 62327 15845
rect 72744 13884 72808 15862
rect 81526 13892 81593 15969
rect 9866 13030 9941 13767
rect 20298 13056 20365 13769
rect 30790 13058 30857 13795
rect 41310 13064 41377 13797
rect 49945 13795 51839 13862
rect 60411 13797 62327 13864
rect 70826 13820 72818 13884
rect 81405 13825 81593 13892
rect 9866 12966 10716 13030
rect 20298 12989 21193 13056
rect 30790 12995 31620 13058
rect 41310 12997 42169 13064
rect 51772 13058 51839 13795
rect 62262 13084 62326 13797
rect 72754 13086 72818 13820
rect 30857 12994 31620 12995
rect 51772 12991 52605 13058
rect 62262 13020 63078 13084
rect 72754 13022 73556 13086
rect 10399 7814 10466 9890
rect 6703 7747 10466 7814
rect 20875 7782 20942 9892
rect 31372 7854 31439 9918
rect 462 -198 526 5866
rect 6703 3864 6770 7747
rect 17221 7715 20942 7782
rect 27717 7787 31439 7854
rect 41860 7844 41927 9920
rect 52338 7876 52405 9918
rect 6703 3791 6770 3797
rect 1975 1941 1981 2008
rect 2048 1941 2054 2008
rect 10944 -198 11008 5862
rect 17221 3834 17288 7715
rect 17221 3761 17288 3767
rect 12451 1931 12457 1998
rect 12524 1931 12530 1998
rect 21428 -198 21492 5930
rect 27717 3844 27784 7787
rect 38171 7777 41927 7844
rect 48635 7809 52405 7876
rect 62808 7834 62875 9920
rect 27717 3771 27784 3777
rect 22937 1963 22943 2030
rect 23010 1963 23016 2030
rect 31910 -198 31974 5892
rect 38171 3896 38238 7777
rect 38171 3823 38238 3829
rect 33409 2030 33476 2036
rect 33409 1957 33476 1963
rect 42388 -198 42452 5892
rect 48635 3852 48702 7809
rect 59131 7767 62875 7834
rect 73293 7796 73360 9946
rect 83780 7876 83847 9948
rect 48635 3779 48702 3785
rect 43875 1965 43881 2032
rect 43948 1965 43954 2032
rect 52870 -198 52934 5950
rect 59131 3864 59198 7767
rect 69647 7703 73360 7796
rect 80131 7809 83847 7876
rect 59131 3791 59198 3797
rect 54391 1975 54397 2042
rect 54464 1975 54470 2042
rect 63354 -198 63418 5930
rect 69647 3914 69714 7703
rect 69647 3841 69714 3847
rect 64855 2005 64861 2072
rect 64928 2005 64934 2072
rect 73836 -198 73900 5948
rect 80131 3894 80198 7809
rect 80131 3821 80198 3827
rect 75331 1995 75337 2062
rect 75404 1995 75410 2062
rect 462 -262 73900 -198
<< via1 >>
rect 6703 3797 6770 3864
rect 1981 1941 2048 2008
rect 17221 3767 17288 3834
rect 12457 1931 12524 1998
rect 27717 3777 27784 3844
rect 22943 1963 23010 2030
rect 38171 3829 38238 3896
rect 33409 1963 33476 2030
rect 48635 3785 48702 3852
rect 43881 1965 43948 2032
rect 59131 3797 59198 3864
rect 54397 1975 54464 2042
rect 69647 3847 69714 3914
rect 64861 2005 64928 2072
rect 80131 3827 80198 3894
rect 75337 1995 75404 2062
<< metal2 >>
rect 1981 3797 6703 3864
rect 6770 3797 6776 3864
rect 1981 2008 2048 3797
rect 1981 1935 2048 1941
rect 12457 3767 17221 3834
rect 17288 3767 17294 3834
rect 22943 3777 27717 3844
rect 27784 3777 27790 3844
rect 33409 3829 38171 3896
rect 38238 3829 38244 3896
rect 12457 1998 12524 3767
rect 22943 2030 23010 3777
rect 33409 2030 33476 3829
rect 43881 3785 48635 3852
rect 48702 3785 48708 3852
rect 54397 3797 59131 3864
rect 59198 3797 59204 3864
rect 64861 3847 69647 3914
rect 69714 3847 69720 3914
rect 43881 2032 43948 3785
rect 33403 1963 33409 2030
rect 33476 1963 33482 2030
rect 54397 2042 54464 3797
rect 64861 2072 64928 3847
rect 64861 1999 64928 2005
rect 75337 3827 80131 3894
rect 80198 3827 80204 3894
rect 75337 2062 75404 3827
rect 75337 1989 75404 1995
rect 54397 1969 54464 1975
rect 22943 1957 23010 1963
rect 43881 1959 43948 1965
rect 12457 1925 12524 1931
use JNW_GR03_DFLIPFLIP_F_R  JNW_GR03_DFLIPFLIP_F_R_4
timestamp 1744305162
transform 1 0 31446 0 1 11862
box 0 -11832 10481 3926
use JNW_GR03_DFLIPFLIP_F_R  JNW_GR03_DFLIPFLIP_F_R_5
timestamp 1744305162
transform 1 0 20964 0 1 11860
box 0 -11832 10481 3926
use JNW_GR03_DFLIPFLIP_F_R  JNW_GR03_DFLIPFLIP_F_R_6
timestamp 1744305162
transform 1 0 10480 0 1 11834
box 0 -11832 10481 3926
use JNW_GR03_DFLIPFLIP_F_R  JNW_GR03_DFLIPFLIP_F_R_7
timestamp 1744305162
transform 1 0 -2 0 1 11832
box 0 -11832 10481 3926
use JNW_GR03_DFLIPFLIP_F_R  JNW_GR03_DFLIPFLIP_F_R_8
timestamp 1744305162
transform 1 0 41924 0 1 11860
box 0 -11832 10481 3926
use JNW_GR03_DFLIPFLIP_F_R  JNW_GR03_DFLIPFLIP_F_R_9
timestamp 1744305162
transform 1 0 52406 0 1 11862
box 0 -11832 10481 3926
use JNW_GR03_DFLIPFLIP_F_R  JNW_GR03_DFLIPFLIP_F_R_10
timestamp 1744305162
transform 1 0 62890 0 1 11888
box 0 -11832 10481 3926
use JNW_GR03_DFLIPFLIP_F_R  JNW_GR03_DFLIPFLIP_F_R_11
timestamp 1744305162
transform 1 0 73372 0 1 11890
box 0 -11832 10481 3926
<< labels >>
flabel metal1 81526 15902 81593 15969 0 FreeSans 1600 0 0 0 B7
flabel metal1 72744 15798 72808 15862 0 FreeSans 1600 0 0 0 B6
flabel metal1 62260 15778 62327 15845 0 FreeSans 1600 0 0 0 B5
flabel metal1 51772 15768 51839 15835 0 FreeSans 1600 0 0 0 B4
flabel metal1 41310 15768 41377 15835 0 FreeSans 1600 0 0 0 B3
flabel metal1 30790 15778 30857 15845 0 FreeSans 1600 0 0 0 B2
flabel metal1 20298 15698 20365 15765 0 FreeSans 1600 0 0 0 B1
flabel metal1 9866 15712 9941 15787 0 FreeSans 1600 0 0 0 B0
<< end >>
