*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_GR03_DFLIPFLOP_R_R_lpe.spi
#else
.include ../../../work/xsch/JNW_GR03_DFLIPFLOP_R_R.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-3

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD  VSS   dc 1.8
VCLK CLK  0     pulse(0.1 1.7 20n 2n 2n 20n  150n)
VRST RST  0     pulse(0.1 1.7 0   2n 2n 350n 1u)
VD   D    0     pulse(0.1 1.7 0   2n 2n 150n 300n)

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save v(CLK)
.save v(RST)
.save v(D)
.save v(Q)
.save v(NOT_Q)


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 1n 1u 0


tran 2n 2u 1p
write
quit


.endc

.end
