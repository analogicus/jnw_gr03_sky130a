** sch_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_GR03_SKY130A/JNW_GR03_TB.sch
.subckt JNW_GR03_TB VDD VSS I_TEMP
*.ipin VDD
*.ipin VSS
*.opin I_TEMP
x4 GS2 VR1 VSS JNWTR_RPPO4
x5<1> VD1 net1 VDD VDD JNWATR_PCH_4C5F0
x5<0> VD1 net1 VDD VDD JNWATR_PCH_4C5F0
x2<1> VR1 net1 VDD VDD JNWATR_PCH_4C5F0
x2<0> VR1 net1 VDD VDD JNWATR_PCH_4C5F0
x6<1> net1 net1 VDD VDD JNWATR_PCH_4C5F0
x6<0> net1 net1 VDD VDD JNWATR_PCH_4C5F0
x7 net1 net2 VSS VSS JNWATR_NCH_4C5F0
x8 VSS net2 JNWTR_CAPX1
x1<1> I_TEMP net1 VDD VDD JNWATR_PCH_4C5F0
x1<0> I_TEMP net1 VDD VDD JNWATR_PCH_4C5F0
x3<1> VD1 VD1 VSS VSS JNWATR_NCH_4C5F0
x3<0> VD1 VD1 VSS VSS JNWATR_NCH_4C5F0
x11 GS2 GS2 VSS VSS JNWATR_NCH_4C5F0
x9 VDD net2 VR1 VD1 VSS JNW_GR03_AMP
.ends

* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO4.sym # of pins=3
** sym_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sym
** sch_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO4.sch
.subckt JNWTR_RPPO4 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES4
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym # of pins=4
** sym_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sym
** sch_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C5F0.sch
.subckt JNWATR_PCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym # of pins=4
** sym_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sym
** sch_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_ATR_SKY130A/JNWATR_NCH_4C5F0.sch
.subckt JNWATR_NCH_4C5F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=0.94 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_CAPX1.sym # of pins=2
** sym_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sym
** sch_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_CAPX1.sch
.subckt JNWTR_CAPX1 A B
*.iopin A
*.iopin B
XC1 B A sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
.ends


* expanding   symbol:  JNW_GR03_SKY130A/JNW_GR03_AMP.sym # of pins=5
** sym_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_GR03_SKY130A/JNW_GR03_AMP.sym
** sch_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_GR03_SKY130A/JNW_GR03_AMP.sch
.subckt JNW_GR03_AMP VDD Vo Vip Vin VSS
*.ipin Vin
*.ipin Vip
*.opin Vo
*.ipin VSS
*.ipin VDD
x2 net2 Vin net1 net1 JNWATR_PCH_4C1F2
x1 net3 Vip net1 net1 JNWATR_PCH_4C1F2
x3 net3 net3 VSS VSS JNWATR_NCH_4C5F0
x4 net2 net2 VSS VSS JNWATR_NCH_4C5F0
x10 Vo net3 VSS VSS JNWATR_NCH_4C5F0
x8 net4 net2 VSS VSS JNWATR_NCH_4C5F0
x7<1> net4 net4 VDD VDD JNWATR_PCH_4C5F0
x7<0> net4 net4 VDD VDD JNWATR_PCH_4C5F0
x9<1> Vo Vo VDD VDD JNWATR_PCH_4C5F0
x9<0> Vo Vo VDD VDD JNWATR_PCH_4C5F0
x1<1> net7<1> net5<1> VDD VDD JNWATR_PCH_4C5F0
x1<0> net7<0> net5<0> VDD VDD JNWATR_PCH_4C5F0
x5<1> net1 net5<1> VDD VDD JNWATR_PCH_4C5F0
x5<0> net1 net5<0> VDD VDD JNWATR_PCH_4C5F0
x9 VSS net6 VSS JNWTR_RPPO4
x12<0> net6 net7<1> VSS JNWTR_RPPO2
x12<1> net6 net7<0> VSS JNWTR_RPPO2
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES4.sym # of pins=3
** sym_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sym
** sch_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RES4.sch
.subckt JNWTR_RES4 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 INT_1 INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_2 INT_2 INT_1 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_3 P INT_2 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends


* expanding   symbol:  JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym # of pins=4
** sym_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sym
** sch_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_ATR_SKY130A/JNWATR_PCH_4C1F2.sch
.subckt JNWATR_PCH_4C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.22 W=3.2 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RPPO2.sym # of pins=3
** sym_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO2.sym
** sch_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RPPO2.sch
.subckt JNWTR_RPPO2 N P B
*.iopin P
*.iopin N
*.iopin B
XXA1 N P B JNWTR_RES2
.ends


* expanding   symbol:  JNW_TR_SKY130A/JNWTR_RES2.sym # of pins=3
** sym_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sym
** sch_path: /home/toushif/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A/JNWTR_RES2.sch
.subckt JNWTR_RES2 N P B
*.iopin N
*.iopin P
*.iopin B
XR1_0 INT_0 N B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
XR1_1 P INT_0 B sky130_fd_pr__res_high_po W=0.36 L=7.36 mult=1 m=1
.ends

.end
