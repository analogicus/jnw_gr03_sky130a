magic
tech sky130A
magscale 1 2
timestamp 1744292387
<< locali >>
rect 1200 3734 2272 3926
rect 3944 3922 4136 3926
rect 1200 2154 1934 3734
rect 3142 3730 6766 3922
rect 1200 2132 1392 2154
rect 1606 556 1934 2154
rect 3944 2294 4316 3730
rect 3944 2114 3950 2294
rect 4310 2114 4316 2294
rect 3944 2108 4316 2114
rect 2420 1932 6375 1999
rect 1606 376 1612 556
rect 1792 546 1934 556
rect 1606 370 1748 376
rect 1742 366 1748 370
rect 1928 366 1934 546
rect 1742 360 1934 366
rect 1154 4 2296 196
rect 3944 -222 4316 1636
rect 6308 -30 6375 1932
rect 5750 -222 6732 -30
rect 1606 -3984 1934 -362
rect 6308 -2093 6375 -222
rect 6308 -2148 6314 -2093
rect 6369 -2148 6375 -2093
rect 6308 -2153 6375 -2148
rect 5716 -3932 6744 -3740
rect 1336 -4176 2352 -3984
rect 5682 -4166 6112 -3974
rect 5920 -5342 6112 -4166
rect 5760 -5534 6630 -5342
rect 1324 -6304 2284 -6112
rect 1720 -11540 1912 -6304
rect 6438 -7918 6630 -5534
rect 5738 -8110 6630 -7918
rect 1720 -11732 2306 -11540
<< viali >>
rect 3950 2114 4310 2294
rect 2365 1932 2420 1999
rect 1612 546 1792 556
rect 1612 376 1928 546
rect 1748 366 1928 376
rect 3944 1636 4316 1816
rect 1606 -362 1934 -182
rect 6314 -2148 6369 -2093
<< metal1 >>
rect 3944 2294 4316 2306
rect 3944 2114 3950 2294
rect 4310 2114 4316 2294
rect 2359 1999 2426 2011
rect 2359 1932 2365 1999
rect 2420 1932 2426 1999
rect 2359 1920 2426 1932
rect 3121 1927 3587 1994
rect 1360 1133 1916 1196
rect 1674 1132 1916 1133
rect 1980 1132 1986 1196
rect 2373 837 2440 843
rect 2373 764 2440 770
rect 1606 558 1798 568
rect 1606 556 1934 558
rect 1606 376 1612 556
rect 1792 546 1934 556
rect 1606 366 1748 376
rect 1928 366 1934 546
rect 1606 -176 1934 366
rect 3520 118 3587 1927
rect 3944 1822 4316 2114
rect 7562 1935 8209 2002
rect 3932 1816 4328 1822
rect 3932 1636 3944 1816
rect 4316 1636 4328 1816
rect 3932 1630 4328 1636
rect 6790 1219 6857 1225
rect 6790 1146 6857 1152
rect 6032 837 6099 843
rect 3514 51 3520 118
rect 3587 51 3593 118
rect 1594 -182 1946 -176
rect 1594 -362 1606 -182
rect 1934 -362 1946 -182
rect 1594 -368 1946 -362
rect 2367 -1221 2373 -1154
rect 2440 -1221 2446 -1154
rect 6032 -1950 6099 770
rect 6784 414 6857 420
rect 6784 335 6857 341
rect 7932 130 7999 1935
rect 7932 57 7999 63
rect 9864 -424 9936 -418
rect 9864 -1206 9936 -496
rect 6787 -1275 6793 -1208
rect 6860 -1275 6866 -1208
rect 1780 -2026 2231 -1963
rect 5601 -2017 6101 -1950
rect 6162 -2000 6659 -1933
rect 1780 -4049 1843 -2026
rect 1780 -4112 2082 -4049
rect 2145 -4112 2151 -4049
rect 1780 -5112 1843 -4112
rect 1446 -5175 1843 -5112
rect 1780 -9476 1843 -5175
rect 2375 -5186 2442 -5180
rect 6032 -5186 6099 -2017
rect 6026 -5253 6032 -5186
rect 6099 -5253 6105 -5186
rect 2375 -5259 2442 -5253
rect 6162 -5894 6229 -2000
rect 10046 -2009 10481 -1942
rect 1920 -5900 1984 -5894
rect 1984 -5964 2234 -5900
rect 5619 -5961 6229 -5894
rect 6308 -2093 6375 -2081
rect 6308 -2148 6314 -2093
rect 6369 -2148 6375 -2093
rect 1920 -5970 1984 -5964
rect 4870 -7432 4934 -7426
rect 4870 -7546 4934 -7496
rect 2369 -9110 2436 -9104
rect 2369 -9183 2436 -9177
rect 6032 -9110 6099 -5961
rect 6032 -9183 6099 -9177
rect 6308 -7432 6375 -2148
rect 6372 -7496 6375 -7432
rect 1770 -9545 1776 -9476
rect 1845 -9545 1851 -9476
rect 1780 -9661 1843 -9545
rect 1032 -9898 2236 -9834
rect 6308 -9838 6375 -7496
rect 5640 -9905 6375 -9838
<< via1 >>
rect 1916 1132 1980 1196
rect 2373 770 2440 837
rect 6790 1152 6857 1219
rect 6032 770 6099 837
rect 3520 51 3587 118
rect 2373 -1221 2440 -1154
rect 6784 341 6857 414
rect 7932 63 7999 130
rect 9864 -496 9936 -424
rect 6793 -1275 6860 -1208
rect 2082 -4112 2145 -4049
rect 2375 -5253 2442 -5186
rect 6032 -5253 6099 -5186
rect 1920 -5964 1984 -5900
rect 4870 -7496 4934 -7432
rect 2369 -9177 2436 -9110
rect 6032 -9177 6099 -9110
rect 6308 -7496 6372 -7432
rect 1776 -9545 1845 -9476
<< metal2 >>
rect 1916 1196 1980 1202
rect 1916 -2234 1980 1132
rect 6032 1152 6790 1219
rect 6857 1152 6863 1219
rect 6032 837 6099 1152
rect 2367 770 2373 837
rect 2440 770 6032 837
rect 6099 770 6105 837
rect 6778 341 6784 414
rect 6857 341 9937 414
rect 3520 118 3587 124
rect 2373 51 3520 118
rect 2373 -1154 2440 51
rect 3520 45 3587 51
rect 6793 63 7932 130
rect 7999 63 8005 130
rect 2373 -1227 2440 -1221
rect 6793 -1208 6860 63
rect 9864 -424 9937 341
rect 9858 -496 9864 -424
rect 9936 -496 9942 -424
rect 6793 -1281 6860 -1275
rect 1916 -2298 2352 -2234
rect 6384 -2292 6809 -2229
rect 1920 -5900 1984 -2298
rect 2082 -4049 2145 -4043
rect 6384 -4049 6447 -2292
rect 2145 -4112 6447 -4049
rect 2082 -4118 2145 -4112
rect 6032 -5186 6099 -5180
rect 2369 -5253 2375 -5186
rect 2442 -5253 6032 -5186
rect 6032 -5259 6099 -5253
rect 1914 -5964 1920 -5900
rect 1984 -5964 1990 -5900
rect 4864 -7496 4870 -7432
rect 4934 -7496 6308 -7432
rect 6372 -7496 6378 -7432
rect 2363 -9177 2369 -9110
rect 2436 -9177 6032 -9110
rect 6099 -9177 6105 -9110
rect 1776 -9476 1845 -9470
rect 1776 -10122 1845 -9545
rect 1776 -10186 2502 -10122
rect 1776 -10191 2333 -10186
use JNW_GR03_NAND3  JNW_GR03_NAND3_0
timestamp 1744292387
transform 1 0 2028 0 1 -11832
box -2 0 4018 3914
use JNW_GR03_NAND3  JNW_GR03_NAND3_1
timestamp 1744292387
transform 1 0 6450 0 1 -3936
box -2 0 4018 3914
use JNW_GR03_NAND3  JNW_GR03_NAND3_2
timestamp 1744292387
transform 1 0 2028 0 1 -7888
box -2 0 4018 3914
use JNW_GR03_NAND3  JNW_GR03_NAND3_3
timestamp 1744292387
transform 1 0 2028 0 1 -3944
box -2 0 4018 3914
use JNW_GR03_NAND  JNW_GR03_NAND_0
timestamp 1744289480
transform 1 0 6634 0 1 1038
box -186 -1030 1334 2884
use JNW_GR03_NAND  JNW_GR03_NAND_1
timestamp 1744289480
transform 1 0 2212 0 1 1030
box -186 -1030 1334 2884
use JNW_GR03_NOT  JNW_GR03_NOT_0
timestamp 1744287221
transform 1 0 120 0 1 -5148
box 0 -1160 1520 1164
use JNW_GR03_NOT  JNW_GR03_NOT_1
timestamp 1744287221
transform 1 0 0 0 1 1160
box 0 -1160 1520 1164
<< labels >>
flabel space 94 1132 158 1196 0 FreeSans 1600 0 0 0 CLK
flabel metal1 1032 -9898 1096 -9834 0 FreeSans 1600 0 0 0 D
flabel space 222 -5176 286 -5112 0 FreeSans 1600 0 0 0 RST
flabel metal1 8142 1935 8209 2002 0 FreeSans 1600 0 0 0 Q
flabel metal1 10414 -2009 10481 -1942 0 FreeSans 1600 0 0 0 NOT_Q
<< end >>
