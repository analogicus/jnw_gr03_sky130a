magic
tech sky130A
magscale 1 2
timestamp 1744318479
<< locali >>
rect -1562 6568 4844 6648
rect -1562 6388 -1024 6568
rect -844 6552 4844 6568
rect -844 6546 3786 6552
rect -844 6388 2536 6546
rect -1562 6366 2536 6388
rect 2716 6372 3786 6546
rect 3966 6372 4844 6552
rect 2716 6366 4844 6372
rect -1562 6328 4844 6366
rect -1414 5790 -1222 6328
rect -262 5838 -70 6328
rect 2146 6036 2338 6328
rect 3298 5988 3588 6328
rect 4548 6000 4740 6328
rect 360 4240 552 4584
rect 1512 4240 1704 4598
rect 356 4048 1704 4240
rect 2146 3500 2338 3704
rect 3298 3500 3590 3734
rect 4550 3500 4742 3686
rect 2146 3320 2536 3500
rect 2716 3496 4742 3500
rect 2716 3320 3788 3496
rect 2146 3316 3788 3320
rect 3968 3316 4742 3496
rect 2146 3314 4742 3316
rect 2148 3308 4742 3314
rect 4344 3130 4554 3308
rect 4344 2950 4370 3130
rect 4550 2950 4554 3130
rect 4344 105 4554 2950
rect -1527 -105 4587 105
<< viali >>
rect -1024 6388 -844 6568
rect 2536 6366 2716 6546
rect 3786 6372 3966 6552
rect 380 5327 531 5478
rect 2536 3320 2716 3500
rect 3788 3316 3968 3496
rect -1102 2962 -922 3142
rect -638 2950 -458 3130
rect 422 2950 602 3130
rect 3892 2950 4072 3130
rect 4370 2950 4550 3130
<< metal1 >>
rect -1030 6568 -838 6580
rect -1030 6388 -1024 6568
rect -844 6388 -838 6568
rect -1030 5624 -838 6388
rect 2530 6546 2722 6558
rect 2530 6366 2536 6546
rect 2716 6366 2722 6546
rect 1140 5934 1309 5940
rect -1158 5008 -1094 5404
rect -1030 4760 -838 5548
rect -631 5484 -468 5914
rect 626 5890 678 5896
rect 626 5832 678 5838
rect 2530 5820 2722 6366
rect 3780 6552 3972 6564
rect 3780 6372 3786 6552
rect 3966 6372 3972 6552
rect 3780 5784 3972 6372
rect -631 5315 -468 5321
rect 374 5484 537 5490
rect 760 5484 923 5490
rect 374 5315 537 5321
rect 746 5321 760 5396
rect 923 5321 936 5396
rect 746 5062 936 5321
rect 1140 5292 1309 5765
rect 2402 5298 2466 5532
rect 2914 5298 3106 5698
rect 3652 5298 3716 5564
rect 2402 5234 3716 5298
rect 4164 5298 4356 5714
rect 4164 5234 4790 5298
rect 1137 5179 1312 5185
rect -1158 4210 -1094 4576
rect -1030 4002 -838 4696
rect -1157 3723 -1095 3841
rect -1158 3504 -1094 3712
rect -646 3504 -454 5058
rect 746 4970 914 5062
rect 1137 4873 1312 5004
rect 2914 4790 3106 5234
rect 4164 4822 4356 5234
rect 622 4552 674 4558
rect 622 4494 674 4500
rect 2402 4168 2466 4556
rect 2402 3802 2466 3808
rect 2402 3578 2466 3738
rect -1158 3314 -454 3504
rect -1108 3312 -454 3314
rect 2530 3500 2722 4696
rect 3652 4294 3716 4504
rect 3652 4198 3718 4294
rect 3654 4188 3718 4198
rect 3654 4118 3718 4124
rect 2924 3852 3099 3858
rect 2924 3671 3099 3677
rect 2530 3320 2536 3500
rect 2716 3320 2722 3500
rect -1108 3142 -916 3312
rect 2530 3308 2722 3320
rect 3782 3496 3974 4648
rect 4179 4239 4348 4245
rect 4179 4064 4348 4070
rect 3782 3316 3788 3496
rect 3968 3316 3974 3496
rect 3782 3304 3974 3316
rect -1108 2962 -1102 3142
rect -922 2962 -916 3142
rect 3886 3136 4078 3142
rect -1108 2950 -916 2962
rect -650 3130 626 3136
rect -650 2950 -638 3130
rect -458 2950 422 3130
rect 602 2950 626 3130
rect -650 2944 626 2950
rect 3884 3130 4562 3136
rect 3884 2950 3892 3130
rect 4072 2950 4370 3130
rect 4550 2950 4562 3130
rect 3884 2944 4562 2950
rect 3886 2938 4078 2944
<< via1 >>
rect 626 5838 678 5890
rect 1140 5765 1309 5934
rect -631 5321 -468 5484
rect 374 5478 537 5484
rect 374 5327 380 5478
rect 380 5327 531 5478
rect 531 5327 537 5478
rect 374 5321 537 5327
rect 760 5321 923 5484
rect 1137 5004 1312 5179
rect 622 4500 674 4552
rect 2402 3738 2466 3802
rect 3654 4124 3718 4188
rect 2924 3677 3099 3852
rect 4179 4070 4348 4239
<< metal2 >>
rect 620 5886 626 5890
rect -1484 5842 626 5886
rect 620 5838 626 5842
rect 678 5838 684 5890
rect 1134 5765 1140 5934
rect 1309 5765 2000 5934
rect -637 5321 -631 5484
rect -468 5321 374 5484
rect 537 5321 760 5484
rect 923 5321 929 5484
rect 1131 5004 1137 5179
rect 1312 5004 1665 5179
rect 616 4548 622 4552
rect -1518 4503 622 4548
rect 616 4500 622 4503
rect 674 4500 680 4552
rect 1490 3852 1665 5004
rect 1831 4239 2000 5765
rect 1831 4188 4179 4239
rect 1831 4124 3654 4188
rect 3718 4124 4179 4188
rect 1831 4070 4179 4124
rect 4348 4070 4354 4239
rect 1490 3802 2924 3852
rect 1490 3738 2402 3802
rect 2466 3738 2924 3802
rect 1490 3677 2924 3738
rect 3099 3677 3105 3852
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1737385461
transform 1 0 2242 0 1 3534
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1 ../JNW_ATR_SKY130A
timestamp 1737385461
transform 1 0 2242 0 1 4332
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2 ../JNW_ATR_SKY130A
timestamp 1737385461
transform 1 0 3494 0 1 3534
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3 ../JNW_ATR_SKY130A
timestamp 1737385461
transform 1 0 3492 0 1 4332
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  JNWATR_PCH_4C1F2_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 456 0 1 4432
box -184 -128 1336 928
use JNWATR_PCH_4C1F2  JNWATR_PCH_4C1F2_1 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 456 0 1 5188
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1318 0 1 3594
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_1 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1318 0 1 5190
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_2 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1318 0 1 4392
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_3 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 3492 0 1 5388
box -184 -128 1336 928
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_4 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 2242 0 1 5388
box -184 -128 1336 928
use JNWTR_RPPO2  JNWTR_RPPO2_0 ../JNW_TR_SKY130A
timestamp 1744275334
transform -1 0 -54 0 1 0
box 0 0 1448 3440
use JNWTR_RPPO16  JNWTR_RPPO16_0 ../JNW_TR_SKY130A
timestamp 1744275334
transform -1 0 4472 0 1 0
box 0 0 4472 3440
<< labels >>
flabel metal2 -1484 5842 -1440 5886 0 FreeSans 1600 0 0 0 Vip
flabel metal2 -1513 4503 -1463 4548 0 FreeSans 1600 0 0 0 Vin
flabel locali -1562 6328 -1242 6648 0 FreeSans 1600 0 0 0 VDD
flabel locali -1527 -105 -1317 105 0 FreeSans 1600 0 0 0 VSS
<< end >>
