magic
tech sky130A
magscale 1 2
timestamp 1744289412
<< metal1 >>
rect 1079 1927 1657 1994
rect 2175 1993 2459 2002
rect 2175 1928 2381 1993
rect 2446 1928 2459 1993
rect 2175 1919 2459 1928
rect 2644 1710 2708 2044
rect 2837 1993 2902 1999
rect 2837 1922 2902 1928
rect 2644 1640 2708 1646
<< via1 >>
rect 2381 1928 2446 1993
rect 2837 1928 2902 1993
rect 2644 1646 2708 1710
<< metal2 >>
rect 2381 1993 2446 1999
rect 2446 1928 2837 1993
rect 2902 1928 2908 1993
rect 2381 1922 2446 1928
rect 234 1646 2644 1710
rect 2708 1646 2714 1710
use JNW_GR03_NAND  JNW_GR03_NAND_0
timestamp 1744288710
transform 1 0 2684 0 1 1030
box -186 -1030 1334 2884
use JNW_GR03_NAND  JNW_GR03_NAND_1
timestamp 1744288710
transform 1 0 184 0 1 1030
box -186 -1030 1334 2884
use JNW_GR03_NAND  JNW_GR03_NAND_2
timestamp 1744288710
transform 1 0 1434 0 1 1030
box -186 -1030 1334 2884
<< labels >>
flabel metal2 234 1646 298 1710 0 FreeSans 1600 0 0 0 C
flabel space 144 1942 208 2006 0 FreeSans 1600 0 0 0 B
flabel space 342 2768 406 2832 0 FreeSans 1600 0 0 0 A
<< end >>
