magic
tech sky130A
magscale 1 2
timestamp 1744548282
<< locali >>
rect 88 9282 4160 9474
rect 88 9122 280 9282
rect 88 6508 280 7032
rect 1112 6540 1304 7068
rect 1476 6530 1668 7036
rect 2500 6530 2692 7048
rect 2868 6534 3060 7032
rect 3892 6514 4084 7068
rect -1432 5594 -1240 6072
rect -1505 194 645 204
rect -1505 14 -1042 194
rect -862 14 645 194
rect -1505 -6 645 14
<< viali >>
rect -2422 8922 -2242 9102
rect -688 8912 -508 9092
rect 1866 6524 2046 6704
rect 3258 6536 3438 6716
rect 5963 591 6069 697
rect -1042 14 -862 194
<< metal1 >>
rect -2428 9102 -2236 9114
rect -2428 8922 -2422 9102
rect -2242 8922 -2236 9102
rect -2428 6324 -2236 8922
rect -694 9098 -502 9104
rect 722 8906 728 9098
rect 920 8906 926 9098
rect -694 8900 -502 8906
rect 344 6982 408 8694
rect 348 6978 404 6982
rect 348 6916 404 6922
rect 472 6486 664 8852
rect 728 7410 920 8810
rect 1732 6978 1796 8668
rect 1732 6950 1736 6978
rect 1792 6950 1796 6978
rect 1736 6916 1792 6922
rect 1860 6704 2052 9062
rect 2116 7330 2308 8810
rect 3124 7512 3188 8670
rect 1860 6524 1866 6704
rect 2046 6524 2052 6704
rect 1860 6512 2052 6524
rect 2192 6340 2256 7134
rect 3124 6978 3180 6984
rect 3252 6978 3444 8794
rect 3508 7342 3700 8832
rect 3124 6916 3180 6922
rect 3252 6716 3444 6922
rect 3252 6536 3258 6716
rect 3438 6536 3444 6716
rect 3252 6524 3444 6536
rect -2428 6132 -472 6324
rect -1176 5622 -1112 6132
rect -664 5466 -472 6132
rect 1668 6276 2256 6340
rect -1176 4758 -1112 5242
rect -1048 4721 -856 5114
rect -664 4721 -472 5302
rect -491 4529 -472 4721
rect 1668 4638 1732 6276
rect 5816 6110 5822 6166
rect 5878 6110 5884 6166
rect 6130 5393 6141 5397
rect 6130 5333 6131 5393
rect 6147 5302 6163 5421
rect 6266 5302 6272 5421
rect 2178 4638 2242 4724
rect 1668 4574 2242 4638
rect -1176 1190 -1112 4322
rect -1175 833 -1123 839
rect -1175 775 -1123 781
rect -1048 194 -856 4529
rect -664 1312 -472 4529
rect 5951 911 5957 1029
rect 6075 911 6081 1029
rect -587 781 -581 833
rect -529 781 -523 833
rect 5957 697 6075 911
rect 5957 591 5963 697
rect 6069 591 6075 697
rect 5957 579 6075 591
rect -1048 14 -1042 194
rect -862 14 -856 194
rect -1048 2 -856 14
<< via1 >>
rect -694 9092 -502 9098
rect -694 8912 -688 9092
rect -688 8912 -508 9092
rect -508 8912 -502 9092
rect -694 8906 -502 8912
rect 728 8906 920 9098
rect 348 6922 404 6978
rect 1736 6922 1792 6978
rect 3124 6922 3180 6978
rect 5822 6110 5878 6166
rect 6163 5302 6266 5421
rect -1175 781 -1123 833
rect 5957 911 6075 1029
rect -581 781 -529 833
<< metal2 >>
rect 728 9098 920 9104
rect -700 8906 -694 9098
rect -502 8906 728 9098
rect -206 6064 -14 8906
rect 728 8900 920 8906
rect 342 6922 348 6978
rect 404 6922 1736 6978
rect 1792 6922 3124 6978
rect 3180 6922 5896 6978
rect 5822 6166 5878 6922
rect 5822 6104 5878 6110
rect -210 5985 -14 6064
rect -210 5941 362 5985
rect -210 5872 -14 5941
rect 6163 5421 6266 5427
rect 6163 5238 6266 5302
rect 6163 5136 6266 5145
rect -266 4602 328 4647
rect -581 833 -529 839
rect -1181 781 -1175 833
rect -1123 829 -1117 833
rect -1123 784 -581 829
rect -1123 781 -1117 784
rect -266 829 -221 4602
rect 5957 1354 6075 1359
rect 5953 1246 5962 1354
rect 6070 1246 6079 1354
rect 5957 1029 6075 1246
rect 5957 905 6075 911
rect -529 784 -221 829
rect -581 775 -529 781
<< via2 >>
rect 6163 5145 6266 5238
rect 5962 1246 6070 1354
<< metal3 >>
rect 6158 5238 6271 5243
rect 6158 5145 6163 5238
rect 6266 5145 6271 5238
rect 6158 5140 6271 5145
rect 6163 3057 6266 5140
rect 4655 2871 6266 3057
rect 6163 2701 6266 2871
rect 5957 1696 6075 1697
rect 5952 1580 5958 1696
rect 6074 1580 6080 1696
rect 5957 1354 6075 1580
rect 5957 1246 5962 1354
rect 6070 1246 6075 1354
rect 5957 1241 6075 1246
<< via3 >>
rect 5958 1580 6074 1696
<< metal4 >>
rect 4932 1978 6075 2096
rect 5957 1696 6075 1978
rect 5957 1580 5958 1696
rect 6074 1580 6075 1696
rect 5957 1579 6075 1580
use JNW_GR03_AMP  JNW_GR03_AMP_0 ../JNW_GR03_SKY130A
timestamp 1744548282
transform 1 0 1562 0 1 99
box -1562 -105 4844 6648
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1336 0 1 202
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1336 0 1 2596
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1336 0 1 3394
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1336 0 1 4990
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1336 0 1 1798
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_5 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1336 0 1 1000
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_6 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1336 0 1 4192
box -184 -128 1336 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 2964 0 1 6874
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_1 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 2964 0 1 7676
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_2 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 184 0 1 6874
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_3 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 184 0 1 7676
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_4 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 1572 0 1 6874
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_5 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 1572 0 1 7676
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_6 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 2964 0 1 8474
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_7 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 1572 0 1 8474
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_8 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 184 0 1 8474
box -184 -128 1208 928
use JNWTR_CAPX1  JNWTR_CAPX1_0 ../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 3932 0 1 1976
box 0 0 1080 1080
use JNWTR_CAPX1  JNWTR_CAPX1_1 ../JNW_TR_SKY130A
timestamp 1737500400
transform 1 0 5242 0 1 1978
box 0 0 1080 1080
use JNWTR_RPPO8  JNWTR_RPPO8_0 ../JNW_TR_SKY130A
timestamp 1744548282
transform 1 0 -2836 0 1 5974
box 0 0 2744 3440
<< labels >>
flabel space 3508 8906 3700 9234 0 FreeSans 1600 0 0 0 I_TEMP
<< end >>
