magic
tech sky130A
timestamp 1744272350
<< error_s >>
rect 3969 2593 4045 4153
rect 4736 3213 5496 3336
rect 4640 975 5400 1067
<< locali >>
rect 1337 4093 1697 4242
rect 4393 4105 4489 4108
rect 1337 3973 2091 4093
rect 4393 4015 4396 4105
rect 4486 4015 4489 4105
rect 1337 443 1697 3973
rect 4393 3954 4489 4015
rect 1824 443 1920 2431
rect 1336 371 1920 443
rect 2400 371 2496 2431
rect 1336 370 2496 371
rect 1336 280 2019 370
rect 2109 280 2496 370
rect 1336 275 2496 280
<< viali >>
rect 3724 3973 3838 4093
rect 4196 3976 4310 4090
rect 4396 4015 4486 4105
rect 2019 280 2109 370
<< metal1 >>
rect 4393 4108 4489 4111
rect 3721 4093 3841 4099
rect 3721 3973 3724 4093
rect 3838 4090 4316 4093
rect 3838 3976 4196 4090
rect 4310 3976 4316 4090
rect 4982 4012 4985 4108
rect 5081 4012 5084 4108
rect 4393 4009 4489 4012
rect 3838 3973 4316 3976
rect 3721 3967 3841 3973
rect 2016 370 2112 2171
rect 2016 280 2019 370
rect 2109 280 2112 370
rect 2016 274 2112 280
<< via1 >>
rect 4393 4105 4489 4108
rect 4393 4015 4396 4105
rect 4396 4015 4486 4105
rect 4486 4015 4489 4105
rect 4393 4012 4489 4015
rect 4985 4012 5081 4108
<< metal2 >>
rect 4985 4108 5081 4111
rect 4390 4012 4393 4108
rect 4489 4012 4985 4108
rect 4985 4009 5081 4012
use JNWATR_PCH_4C5F0  JNWATR_PCH_4C5F0_0 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 5033 0 1 4821
box -92 -64 668 464
use JNWATR_PCH_4C1F2  x1 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 4710 0 1 476
box -92 -64 668 464
use JNWATR_PCH_4C1F2  x2
timestamp 1734044400
transform 1 0 4732 0 1 1039
box -92 -64 668 464
use JNWATR_NCH_4C5F0  x3 ../JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 1872 0 1 912
box -92 -64 668 464
use JNWATR_NCH_4C5F0  x4
timestamp 1734044400
transform 1 0 1872 0 1 1477
box -92 -64 668 464
use JNWATR_PCH_4C5F0  x5[0:0]
timestamp 1734044400
transform 1 0 4824 0 1 2217
box -92 -64 668 464
use JNWATR_NCH_4C5F0  x6
timestamp 1734044400
transform 1 0 1872 0 1 393
box -92 -64 668 464
use JNWATR_PCH_4C5F0  x7[0:0]
timestamp 1734044400
transform 1 0 4824 0 1 2745
box -92 -64 668 464
use JNWATR_PCH_4C5F0  x8[0:0]
timestamp 1734044400
transform 1 0 4828 0 1 3277
box -92 -64 668 464
use JNWATR_NCH_4C5F0  x8
timestamp 1734044400
transform 1 0 1872 0 1 2011
box -92 -64 668 464
use JNWATR_PCH_4C5F0  x9[1:0]
timestamp 1734044400
transform 1 0 4841 0 1 3764
box -92 -64 668 464
use JNWTR_RPPO2  x11 ../JNW_TR_SKY130A
timestamp 1743080447
transform 1 0 3989 0 1 2513
box 0 0 724 1720
use JNWTR_RPPO16  x12 ../JNW_TR_SKY130A
timestamp 1743080447
transform 1 0 1789 0 1 2513
box 0 0 2236 1720
<< properties >>
string FIXED_BBOX 0 0 7568 1720
<< end >>
