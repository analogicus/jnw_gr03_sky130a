magic
tech sky130A
magscale 1 2
timestamp 1744320150
<< locali >>
rect 88 9282 4160 9474
rect 88 9122 280 9282
rect 88 6508 280 7032
rect 1112 6540 1304 7068
rect 1476 6530 1668 7036
rect 2500 6530 2692 7048
rect 2868 6534 3060 7032
rect 3892 6514 4084 7068
rect -1432 5594 -1240 6072
rect -1505 -6 645 204
<< viali >>
rect -2422 8922 -2242 9102
rect -688 8912 -508 9092
rect 1866 6524 2046 6704
rect 3258 6536 3438 6716
<< metal1 >>
rect -2428 9102 -2236 9114
rect -2428 8922 -2422 9102
rect -2242 8922 -2236 9102
rect -2428 6324 -2236 8922
rect -694 9098 -502 9104
rect 722 8906 728 9098
rect 920 8906 926 9098
rect -694 8900 -502 8906
rect 344 6982 408 8694
rect 348 6978 404 6982
rect 348 6916 404 6922
rect 472 6486 664 8852
rect 728 7410 920 8810
rect 1732 6978 1796 8668
rect 1732 6950 1736 6978
rect 1792 6950 1796 6978
rect 1736 6916 1792 6922
rect 1860 6704 2052 9062
rect 2116 7330 2308 8810
rect 3124 6978 3180 6984
rect 3252 6978 3444 8794
rect 3508 7342 3700 8832
rect 3124 6916 3180 6922
rect 1860 6524 1866 6704
rect 2046 6524 2052 6704
rect 3252 6716 3444 6922
rect 3252 6536 3258 6716
rect 3438 6536 3444 6716
rect 3252 6524 3444 6536
rect 1860 6512 2052 6524
rect -2428 6132 -856 6324
rect -1176 5740 -1112 5746
rect -1176 5670 -1112 5676
rect -1048 5444 -856 6132
rect 5816 6110 5822 6166
rect 5878 6110 5884 6166
rect -672 5536 -666 5728
rect -474 5536 -468 5728
rect -1171 4652 -1119 4658
rect -1171 4594 -1119 4600
rect -1176 796 -1112 4322
rect -1048 12 -856 5354
rect -664 4651 -472 4846
rect -664 4599 -613 4651
rect -561 4599 -472 4651
rect -664 712 -472 4599
<< via1 >>
rect -694 9092 -502 9098
rect -694 8912 -688 9092
rect -688 8912 -508 9092
rect -508 8912 -502 9092
rect -694 8906 -502 8912
rect 728 8906 920 9098
rect 348 6922 404 6978
rect 1736 6922 1792 6978
rect 3124 6922 3180 6978
rect -1176 5676 -1112 5740
rect 5822 6110 5878 6166
rect -666 5536 -474 5728
rect -1171 4600 -1119 4652
rect -613 4599 -561 4651
<< metal2 >>
rect 728 9098 920 9104
rect -700 8906 -694 9098
rect -502 8906 728 9098
rect -206 6064 -14 8906
rect 728 8900 920 8906
rect 342 6922 348 6978
rect 404 6922 1736 6978
rect 1792 6922 3124 6978
rect 3180 6922 5896 6978
rect 5822 6166 5878 6922
rect 5822 6104 5878 6110
rect -666 5985 -14 6064
rect -666 5968 362 5985
rect -1176 5941 362 5968
rect -1176 5904 -14 5941
rect -1176 5740 -1112 5904
rect -666 5872 -14 5904
rect -1182 5676 -1176 5740
rect -1112 5676 -1106 5740
rect -666 5728 -474 5872
rect -666 5530 -474 5536
rect -1177 4600 -1171 4652
rect -1119 4648 -1113 4652
rect -619 4648 -613 4651
rect -1119 4603 -613 4648
rect -1119 4600 -1113 4603
rect -619 4599 -613 4603
rect -561 4647 -555 4651
rect -561 4602 328 4647
rect -561 4599 -555 4602
use JNW_GR03_AMP  JNW_GR03_AMP_0
timestamp 1744318479
transform 1 0 1562 0 1 99
box -1562 -105 4844 6648
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ~/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_ATR_SKY130A
timestamp 1737385461
transform 1 0 -1336 0 1 202
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_1
timestamp 1737385461
transform 1 0 -1336 0 1 2596
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_2
timestamp 1737385461
transform 1 0 -1336 0 1 3394
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_3
timestamp 1737385461
transform 1 0 -1336 0 1 4990
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_4
timestamp 1737385461
transform 1 0 -1336 0 1 1798
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_5
timestamp 1737385461
transform 1 0 -1336 0 1 1000
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_6
timestamp 1737385461
transform 1 0 -1336 0 1 4192
box -184 -128 1336 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_0 ~/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 2964 0 1 6874
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_1
timestamp 1734044400
transform 1 0 2964 0 1 7676
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_2
timestamp 1734044400
transform 1 0 184 0 1 6874
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_3
timestamp 1734044400
transform 1 0 184 0 1 7676
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_4
timestamp 1734044400
transform 1 0 1572 0 1 6874
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_5
timestamp 1734044400
transform 1 0 1572 0 1 7676
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_6
timestamp 1734044400
transform 1 0 2964 0 1 8474
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_7
timestamp 1734044400
transform 1 0 1572 0 1 8474
box -184 -128 1208 928
use JNWATR_PCH_2C5F0  JNWATR_PCH_2C5F0_8
timestamp 1734044400
transform 1 0 184 0 1 8474
box -184 -128 1208 928
use JNWTR_RPPO8  JNWTR_RPPO8_0 ~/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A
timestamp 1744320150
transform 1 0 -2836 0 1 5974
box 0 0 2744 3440
<< labels >>
flabel space 3508 8906 3700 9234 0 FreeSans 1600 0 0 0 I_TEMP
<< end >>
