magic
tech sky130A
magscale 1 2
timestamp 1744292387
<< metal1 >>
rect 8058 13767 10403 13834
rect 18564 13773 19601 13840
rect 10336 13034 10403 13767
rect 10336 12967 10695 13034
rect 10336 12963 10403 12967
rect 10317 9823 10551 9890
rect 20815 9829 21069 9896
rect 10484 7464 10551 9823
rect 6565 7397 10551 7464
rect -140 6656 398 6720
rect 98 4054 162 6656
rect 98 3990 1452 4054
rect 1516 3990 1522 4054
rect 6565 3842 6632 7397
rect 10038 6658 10886 6722
rect 6804 4054 6868 4060
rect 10038 4054 10102 6658
rect 6868 3990 10102 4054
rect 21002 3990 21069 9829
rect 6804 3984 6868 3990
rect 17259 3923 17265 3990
rect 17332 3923 21069 3990
rect 6565 3769 6632 3775
rect 1315 1927 1321 1994
rect 1388 1927 1394 1994
rect 11679 1951 11685 2018
rect 11752 1951 11758 2018
<< via1 >>
rect 1452 3990 1516 4054
rect 6804 3990 6868 4054
rect 17265 3923 17332 3990
rect 6565 3775 6632 3842
rect 1321 1927 1388 1994
rect 11685 1951 11752 2018
<< metal2 >>
rect 1452 4054 1516 4060
rect 1516 3990 6804 4054
rect 6868 3990 6874 4054
rect 17265 3990 17332 3996
rect 1452 3984 1516 3990
rect 11685 3923 17265 3990
rect 1321 3775 6565 3842
rect 6632 3775 6638 3842
rect 1321 1994 1388 3775
rect 11685 2018 11752 3923
rect 17265 3917 17332 3923
rect 11685 1945 11752 1951
rect 1321 1921 1388 1927
use JNW_GR03_DFLIPFLIP_F_R  JNW_GR03_DFLIPFLIP_F_R_0
timestamp 1744292387
transform 1 0 10502 0 1 11838
box 0 -11832 10481 3926
use JNW_GR03_DFLIPFLIP_F_R  JNW_GR03_DFLIPFLIP_F_R_1
timestamp 1744292387
transform 1 0 0 0 1 11832
box 0 -11832 10481 3926
<< labels >>
flabel metal1 9607 13767 9693 13834 0 FreeSans 1600 0 0 0 B0
flabel metal1 19345 13773 19412 13840 0 FreeSans 1600 0 0 0 B1
<< end >>
