magic
tech sky130A
magscale 1 2
timestamp 1744295509
<< locali >>
rect 2780 5254 3400 5446
rect 1140 3586 1944 3778
rect 1140 2642 1332 3586
rect 894 2450 1332 2642
rect 1140 1562 1612 1754
rect 1420 1502 1612 1562
rect 2768 1536 3346 1728
rect 4248 1536 4846 1728
rect 1420 1310 1996 1502
rect 2844 1310 3432 1502
rect 916 -550 1108 512
rect 916 -742 1954 -550
rect 4654 -614 4846 1536
rect 1762 -2380 1954 -742
rect 4312 -806 4846 -614
rect 2640 -2408 3454 -2216
<< metal1 >>
rect 1476 3454 1888 3518
rect 2788 3459 3030 3526
rect 3097 3459 3103 3526
rect 244 3160 1274 3224
rect 1338 3160 1344 3224
rect 244 2294 308 3160
rect 1476 1744 1540 3454
rect 2026 3224 2090 3230
rect 2026 3154 2090 3160
rect 3218 2454 3282 3592
rect 3414 3526 3481 3532
rect 3414 3453 3481 3459
rect 3992 3176 4056 3182
rect 3992 3106 4056 3112
rect 3218 2384 3282 2390
rect 1470 1680 1476 1744
rect 1540 1680 1546 1744
rect 1226 1451 1695 1514
rect 1476 1310 1540 1316
rect 1476 -416 1540 1246
rect 1632 370 1695 1451
rect 3416 376 3480 382
rect 1632 301 1695 307
rect 2022 370 2085 376
rect 2022 301 2085 307
rect 3416 306 3480 312
rect 3998 -4 4062 2
rect 3998 -74 4062 -68
rect 1214 -480 1884 -416
rect 2788 -485 3283 -418
<< via1 >>
rect 3030 3459 3097 3526
rect 1274 3160 1338 3224
rect 2026 3160 2090 3224
rect 3414 3459 3481 3526
rect 3992 3112 4056 3176
rect 3218 2390 3282 2454
rect 1476 1680 1540 1744
rect 1476 1246 1540 1310
rect 1632 307 1695 370
rect 2022 307 2085 370
rect 3416 312 3480 376
rect 3998 -68 4062 -4
<< metal2 >>
rect 3030 3526 3097 3532
rect 3097 3459 3414 3526
rect 3481 3459 3487 3526
rect 3030 3453 3097 3459
rect 1274 3224 1338 3230
rect 1338 3160 2026 3224
rect 2090 3160 2096 3224
rect 1274 3154 1338 3160
rect 3416 3112 3992 3176
rect 4056 3112 4062 3176
rect 3212 2390 3218 2454
rect 3282 2390 3288 2454
rect 1476 1744 1540 1750
rect 1476 1310 1540 1680
rect 1470 1246 1476 1310
rect 1540 1246 1546 1310
rect 1626 307 1632 370
rect 1695 307 2022 370
rect 2085 307 2091 370
rect 3218 -4 3282 2390
rect 3416 376 3480 3112
rect 3410 312 3416 376
rect 3480 312 3486 376
rect 3218 -68 3998 -4
rect 4062 -68 4068 -4
use JNW_GR03_NAND  JNW_GR03_NAND_0
timestamp 1744289480
transform 1 0 3258 0 1 -1382
box -186 -1030 1334 2884
use JNW_GR03_NAND  JNW_GR03_NAND_1
timestamp 1744289480
transform 1 0 3258 0 1 2562
box -186 -1030 1334 2884
use JNW_GR03_NAND  JNW_GR03_NAND_2
timestamp 1744289480
transform 1 0 1860 0 1 2562
box -186 -1030 1334 2884
use JNW_GR03_NAND  JNW_GR03_NAND_3
timestamp 1744289480
transform 1 0 1860 0 1 -1382
box -186 -1030 1334 2884
use JNW_GR03_NOT  JNW_GR03_NOT_0
timestamp 1744287221
transform 1 0 -100 0 1 1478
box 0 -1160 1520 1164
<< labels >>
flabel metal1 1214 -480 1278 -416 0 FreeSans 1600 0 0 0 E
flabel space -8 1450 56 1514 0 FreeSans 1600 0 0 0 D
flabel space 4171 3459 4248 3526 0 FreeSans 1600 0 0 0 Q
flabel space 4186 -485 4253 -418 0 FreeSans 1600 0 0 0 NOT_Q
<< end >>
