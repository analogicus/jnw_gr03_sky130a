magic
tech sky130A
magscale 1 2
timestamp 1744555364
<< locali >>
rect 2 3713 4806 3802
rect 2 3547 3895 3713
rect 4061 3547 4806 3713
rect 2 3482 4806 3547
rect 4486 3454 4806 3482
rect 4486 3134 10892 3454
rect 4486 2939 7327 3134
rect 10572 2939 10892 3134
rect -1692 2132 -1500 2552
rect -540 2132 -348 2550
rect -1692 2130 -348 2132
rect -1692 1950 -1302 2130
rect -1122 1950 -348 2130
rect -1692 1940 -348 1950
rect -540 740 -348 1940
rect -540 -366 92 740
rect -540 -382 -104 -366
rect -148 -539 -104 -382
rect 69 -539 92 -366
rect -148 -3403 92 -539
rect 4347 -3403 4731 -3284
rect 5890 -3403 6160 21
rect 6528 -3403 7411 -3284
rect 9904 -3403 10664 -3284
rect -148 -3436 10664 -3403
rect -148 -3524 5470 -3436
rect 5558 -3524 10664 -3436
rect -148 -3612 10664 -3524
rect 5 -3613 10664 -3612
<< viali >>
rect 3895 3547 4061 3713
rect 377 2949 568 3128
rect 3895 2953 4061 3131
rect -1302 1950 -1122 2130
rect -104 -539 69 -366
rect 403 -546 576 -361
rect 3895 -527 4061 -361
rect 5470 -3524 5558 -3436
<< metal1 >>
rect 3889 3713 4067 3725
rect 3889 3547 3895 3713
rect 4061 3547 4067 3713
rect 377 3134 568 3151
rect 365 3128 580 3134
rect -1308 2776 -1116 3122
rect -924 3044 -732 3128
rect -924 2944 -866 3044
rect -766 2944 -732 3044
rect -1308 2130 -1116 2712
rect -1308 1950 -1302 2130
rect -1122 1950 -1116 2130
rect -1308 1938 -1116 1950
rect -924 -2366 -732 2944
rect 365 2949 377 3128
rect 568 2949 580 3128
rect 365 2943 580 2949
rect 3889 3131 4067 3547
rect 3889 2953 3895 3131
rect 4061 2953 4067 3131
rect 377 2075 568 2943
rect 3889 2935 4067 2953
rect 377 1899 4067 2075
rect 379 1897 4067 1899
rect 3889 1163 4067 1897
rect 3889 1111 3933 1163
rect 3985 1111 4067 1163
rect 397 -360 582 -349
rect -116 -361 582 -360
rect -116 -366 403 -361
rect -116 -539 -104 -366
rect 69 -539 403 -366
rect -116 -545 403 -539
rect 397 -546 403 -545
rect 576 -546 582 -361
rect 3889 -361 4067 1111
rect 3889 -527 3895 -361
rect 4061 -527 4067 -361
rect 3889 -539 4067 -527
rect 397 -558 582 -546
rect 5464 -3436 5564 -3424
rect 5464 -3524 5470 -3436
rect 5558 -3524 5564 -3436
rect 4866 -3880 4966 -3874
rect 5464 -3880 5564 -3524
rect 4966 -3980 5564 -3880
rect 4866 -3986 4966 -3980
<< via1 >>
rect -866 2944 -766 3044
rect 3933 1111 3985 1163
rect 4866 -3980 4966 -3880
<< metal2 >>
rect -866 3044 -766 3050
rect -866 2537 -766 2944
rect -870 2447 -861 2537
rect -771 2497 -762 2537
rect -771 2453 4612 2497
rect -771 2447 -762 2453
rect -866 2442 -766 2447
rect 3927 1111 3933 1163
rect 3985 1159 3991 1163
rect 3985 1114 4674 1159
rect 3985 1111 3991 1114
rect 4295 -3880 4385 -3876
rect 4290 -3885 4866 -3880
rect 4290 -3975 4295 -3885
rect 4385 -3975 4866 -3885
rect 4290 -3980 4866 -3975
rect 4966 -3980 4972 -3880
rect 4295 -3984 4385 -3980
<< via2 >>
rect -861 2447 -771 2537
rect 4295 -3975 4385 -3885
<< metal3 >>
rect -866 2537 -766 2542
rect -866 2447 -861 2537
rect -771 2447 -766 2537
rect -866 -526 -766 2447
rect 5862 -526 5942 -456
rect 7422 -526 7502 -342
rect 8752 -526 8832 -480
rect 10312 -526 10392 -494
rect -866 -626 10392 -526
rect 5862 -2160 5942 -626
rect 7422 -3394 7502 -626
rect 8752 -3388 8832 -626
rect 10312 -3388 10392 -626
rect 8752 -3394 10707 -3388
rect 3852 -3494 10707 -3394
rect 3761 -3880 3859 -3875
rect 3760 -3881 4390 -3880
rect 3760 -3979 3761 -3881
rect 3859 -3885 4390 -3881
rect 3859 -3975 4295 -3885
rect 4385 -3975 4390 -3885
rect 3859 -3979 4390 -3975
rect 3760 -3980 4390 -3979
rect 3761 -3985 3859 -3980
<< via3 >>
rect 3761 -3979 3859 -3881
<< metal4 >>
rect 5862 -526 5942 -176
rect 7422 -526 7502 -50
rect 8752 -526 8832 -228
rect 10312 -526 10392 -194
rect 5712 -626 10538 -526
rect 5862 -3394 5942 -626
rect 7422 -3394 7502 -626
rect 8752 -3394 8832 -626
rect 10312 -3394 10392 -626
rect 3738 -3494 10754 -3394
rect 3760 -3881 3860 -3494
rect 3760 -3979 3761 -3881
rect 3859 -3979 3860 -3881
rect 3760 -3980 3860 -3979
use JNW_GR03_AMP  JNW_GR03_AMP_0
timestamp 1744555364
transform 1 0 6048 0 1 -3389
box -1562 -105 4844 6648
use JNWATR_NCH_4C5F0  JNWATR_NCH_4C5F0_0 ~/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_ATR_SKY130A
timestamp 1734044400
transform 1 0 -1596 0 1 2368
box -184 -128 1336 928
use JNWTR_CAPX4  JNWTR_CAPX4_0 ~/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A
timestamp 1744555364
transform 1 0 4882 0 1 -3494
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_1
timestamp 1744555364
transform 1 0 7772 0 1 -3494
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_2
timestamp 1744555364
transform 1 0 7764 0 1 -626
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_3
timestamp 1744555364
transform 1 0 1988 0 1 -3494
box 480 0 3120 2640
use JNWTR_CAPX4  JNWTR_CAPX4_4
timestamp 1744555364
transform 1 0 4882 0 1 -626
box 480 0 3120 2640
use JNWTR_RPPO16  JNWTR_RPPO16_0 ~/pro/aicex/ip/jnw_gr03_sky130a/design/JNW_TR_SKY130A
timestamp 1744555364
transform 1 0 -14 0 1 -3494
box 0 0 4472 3440
use JNWTR_RPPO16  JNWTR_RPPO16_1
timestamp 1744555364
transform 1 0 -12 0 1 2
box 0 0 4472 3440
<< labels >>
flabel space -1436 3022 -1372 3086 0 FreeSans 1600 0 0 0 Reset
flabel metal1 -924 2936 -732 3128 0 FreeSans 1600 0 0 0 I_in
<< end >>
