magic
tech sky130A
timestamp 1744283476
<< error_s >>
rect 740 2025 743 2028
rect 737 2022 740 2025
rect 737 1993 740 1996
rect 740 1990 743 1993
rect 1330 1980 1455 2384
rect 1502 2025 1505 2028
rect 1499 2022 1502 2025
rect 1499 1993 1502 1996
rect 1502 1990 1505 1993
rect 2093 1980 2217 2384
rect 2265 2025 2268 2028
rect 2262 2022 2265 2025
rect 2262 1993 2265 1996
rect 2265 1990 2268 1993
rect 568 1856 1328 1980
rect 1330 1856 2090 1980
rect 2093 1856 2853 1980
rect 1330 1325 1455 1853
rect 1502 1380 1505 1383
rect 1499 1377 1502 1380
rect 1499 1348 1502 1351
rect 1502 1345 1505 1348
rect 2093 1325 2217 1853
rect 1375 304 1376 306
rect 2138 304 2139 306
rect 1358 287 1376 289
rect 2121 287 2139 289
<< locali >>
rect 913 2357 2805 2453
rect 615 193 2807 289
<< metal1 >>
rect 1004 1290 1534 1346
rect 1764 1285 2297 1346
<< via1 >>
rect 1502 1348 1534 1380
<< metal2 >>
rect 1534 1348 1727 1380
rect 573 611 941 643
rect 2465 474 2497 646
rect 568 442 2497 474
use JNW_GR03_NAND  x1
timestamp 1744282624
transform 1 0 80 0 1 334
box 488 -144 1250 2119
use JNW_GR03_NAND  x2
timestamp 1744282624
transform 1 0 842 0 1 334
box 488 -144 1250 2119
use JNW_GR03_NAND  x3
timestamp 1744282624
transform 1 0 1605 0 1 334
box 488 -144 1250 2119
<< labels >>
flabel space 2519 1240 2617 1388 0 FreeSans 800 0 0 0 Y
port 1 nsew
flabel locali 948 2362 1210 2452 0 FreeSans 800 0 0 0 VDD
port 2 nsew
flabel space 610 194 782 284 0 FreeSans 800 0 0 0 VSS
port 3 nsew
flabel space 740 1245 771 1380 0 FreeSans 800 0 0 0 A
port 4 nsew
flabel space 571 612 597 641 0 FreeSans 800 0 0 0 B
port 6 nsew
flabel metal2 568 443 597 466 0 FreeSans 800 0 0 0 C
port 7 nsew
<< properties >>
string FIXED_BBOX 0 0 6912 400
<< end >>
